` ifndef _IMEM
` define _IMEM

module IMEM(
		input [7:0] 	IMEM_PC,
		output [31:0]	IMEM_instruction
);

endmodule































	
` endif
